module CSR (
    
);
    
endmodule