//--------------------------- Info ---------------------------//
    //Module Name :　 DMA
    //INFO        :   
    //                
//----------------------- Environment -----------------------//

//------------------------- Module -------------------------//
  module DMA (
    input clk, rst,
    input         DMAEN,
    input         DMASRC,
    input         DMADST,
    input         DMALEN,
    output logic  DMA_interrupt
  );
    
//---------------------- Main code -------------------------//
//-------------------- Slave (CPU2DMA) ---------------------//


//-------------------- Master (CPU2S) ----------------------//
  //--------------------- Arbiter -------------------------//

  endmodule
