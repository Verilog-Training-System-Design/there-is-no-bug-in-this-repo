`ifndef _PARAMETER_SETTING_
`define _PARAMETER_SETTING_

//DATA Parameter
    `define DATA_WIDTH      32
    `define MULT_DATA_WIDTH 64
    `define CSR_REG_WIDTH   64

    `define OP_CODE         7
    `define FUNCTION_3      3
    `define FUNCTION_7      7
    //IEEE 754
    `define EXP             8
    `define FRACTION        23  
    //Memory Define
    `define MEM_ADDR_LEN    14   
`endif
