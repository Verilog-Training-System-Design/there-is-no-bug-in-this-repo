module WDT (
  input     clk,  rst,
  input     clk2, rst2,
  input     WDEN,
  input     WDLIVE,
  input     [31:0]  WTOCNT,
  output    WTO
);
  


  
endmodule